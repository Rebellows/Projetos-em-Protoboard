module dcm (

);

endmodule