module wrapper (
  
);

endmodule