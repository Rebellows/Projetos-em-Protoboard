module dm (
  
);

endmodule